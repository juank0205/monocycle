module mono_tb;

logic clk;
  
endmodule
